// @description
//  ** PART OF **
//  RMR8PM3001A - Taurus 3001
//  (RISC-V 64-bit Privileged Minimal System Processor for T110 ASIC)
//
//  Register Alias Table Global Checkpoints
//
// @author Kumonda221
//

module issue_rat_gc #(
    
) (

);

endmodule
